module sum (
    input data,
    output sum
);
    
endmodule